-------------------------------------------------------------------------------
-- cntr5bit - entity/architecture pair
-------------------------------------------------------------------------------
--  ***************************************************************************
--  ** DISCLAIMER OF LIABILITY                                               **
--  **                                                                       **
--  **  This file contains proprietary and confidential information of       **
--  **  Xilinx, Inc. ("Xilinx"), that is distributed under a license         **
--  **  from Xilinx, and may be used, copied and/or disclosed only           **
--  **  pursuant to the terms of a valid license agreement with Xilinx.      **
--  **                                                                       **
--  **  XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION                **
--  **  ("MATERIALS") "AS IS" WITHOUT WARRANTY OF ANY KIND, EITHER           **
--  **  EXPRESSED, IMPLIED, OR STATUTORY, INCLUDING WITHOUT                  **
--  **  LIMITATION, ANY WARRANTY WITH RESPECT TO NONINFRINGEMENT,            **
--  **  MERCHANTABILITY OR FITNESS FOR ANY PARTICULAR PURPOSE. Xilinx        **
--  **  does not warrant that functions included in the Materials will       **
--  **  meet the requirements of Licensee, or that the operation of the      **
--  **  Materials will be uninterrupted or error-free, or that defects       **
--  **  in the Materials will be corrected. Furthermore, Xilinx does         **
--  **  not warrant or make any representations regarding use, or the        **
--  **  results of the use, of the Materials in terms of correctness,        **
--  **  accuracy, reliability or otherwise.                                  **
--  **                                                                       **
--  **  Xilinx products are not designed or intended to be fail-safe,        **
--  **  or for use in any application requiring fail-safe performance,       **
--  **  such as life-support or safety devices or systems, Class III         **
--  **  medical devices, nuclear facilities, applications related to         **
--  **  the deployment of airbags, or any other applications that could      **
--  **  lead to death, personal injury or severe property or                 **
--  **  environmental damage (individually and collectively, "critical       **
--  **  applications"). Customer assumes the sole risk and liability         **
--  **  of any use of Xilinx products in critical applications,              **
--  **  subject only to applicable laws and regulations governing            **
--  **  limitations on product liability.                                    **
--  **                                                                       **
--  **  Copyright 2010 Xilinx, Inc.                                          **
--  **  All rights reserved.                                                 **
--  **                                                                       **
--  **  This disclaimer and copyright notice must be retained as part        **
--  **  of this file at all times.                                           **
--  ***************************************************************************
--
-------------------------------------------------------------------------------
-- Filename     : cntr5bit.vhd
-- Version      : v2.0
-- 
-- Description  : This file contains the a 5 bit resetable, loadable
--                down counter by 1.
-- VHDL-Standard:   VHDL'93
-------------------------------------------------------------------------------
-- Structure:   
--
--  axi_ethernetlite.vhd
--      \
--      \-- axi_interface.vhd
--      \-- xemac.vhd
--           \
--           \-- mdio_if.vhd
--           \-- emac_dpram.vhd                     
--           \    \                     
--           \    \-- RAMB16_S4_S36
--           \                          
--           \    
--           \-- emac.vhd                     
--                \                     
--                \-- MacAddrRAM                   
--                \-- receive.vhd
--                \      rx_statemachine.vhd
--                \      rx_intrfce.vhd
--                \         async_fifo_fg.vhd
--                \      crcgenrx.vhd
--                \                     
--                \-- transmit.vhd
--                       crcgentx.vhd
--                          crcnibshiftreg
--                       tx_intrfce.vhd
--                          async_fifo_fg.vhd
--                       tx_statemachine.vhd
--                       deferral.vhd
--                          cntr5bit.vhd
--                          defer_state.vhd
--                       bocntr.vhd
--                          lfsr16.vhd
--                       msh_cnt.vhd
--                       ld_arith_reg.vhd
--
-------------------------------------------------------------------------------
-- Author:    PVK
-- History:    
-- PVK        06/07/2010     First Version
-- ^^^^^^
-- First version.  
-- ~~~~~~
-------------------------------------------------------------------------------
-- Naming Conventions:
--      active low signals:                     "*_n"
--      clock signals:                          "Clk", "clk_div#", "clk_#x" 
--      reset signals:                          "Rst", "rst_n" 
--      generics:                               "C_*" 
--      user defined types:                     "*_TYPE" 
--      state machine next state:               "*_ns" 
--      state machine current state:            "*_cs" 
--      combinatorial signals:                  "*_com" 
--      pipelined or register delay signals:    "*_d#" 
--      counter signals:                        "*cnt*"
--      clock enable signals:                   "*_ce" 
--      internal version of output port         "*_i"
--      device pins:                            "*_pin" 
--      ports:                                  - Names begin with Uppercase 
--      processes:                              "*_PROCESS" 
--      component instantiations:               "<ENTITY_>I_<#|FUNC>
-------------------------------------------------------------------------------
-- 
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------------
-- axi_ethernetlite_v3_0_7 library is used for axi_ethernetlite_v3_0_7 
-- component declarations
-------------------------------------------------------------------------------
library axi_ethernetlite_v3_0_7;
use axi_ethernetlite_v3_0_7.mac_pkg.all;

-------------------------------------------------------------------------------
-- Port Declaration
-------------------------------------------------------------------------------
-- Definition of Ports:
--
--  Clk       -- System Clock
--  Rst       -- System Reset
--  Cntout    -- Counter output
--  En        -- Counter enable 
--  Ld        -- Counter load enable
--  Load_in   -- Counter load data
--  Zero      -- Terminal count
-------------------------------------------------------------------------------
-- ENTITY
-------------------------------------------------------------------------------
entity cntr5bit is

  port (
    Clk     : in  std_logic;                  -- input clock
    Rst     : in  std_logic;                  -- reset counter
    Cntout  : out std_logic_vector (0 to 4);
    En      : in  std_logic;                  -- counter down enable by 1
    Ld      : in  std_logic;                  -- load enable
    Load_in : in  std_logic_vector (0 to 4);  -- load input value
    Zero    : out std_logic                  -- terminal count
  );
end cntr5bit;

architecture implementation of cntr5bit is

attribute DowngradeIPIdentifiedWarnings: string;

attribute DowngradeIPIdentifiedWarnings of implementation : architecture is "yes";

-------------------------------------------------------------------------------
--  Constant Declarations
-------------------------------------------------------------------------------
-- Constants used in this design are found in mac_pkg.vhd
-------------------------------------------------------------------------------
-- Signal and Type Declarations
-------------------------------------------------------------------------------
signal count : std_logic_vector(0 to 4);
signal zero_i : std_logic;

begin
Cntout <= count;
 -------------------------------------------------------------------------------
 -- INT_count_PROCESS
 -------------------------------------------------------------------------------
 -- This process assigns the internal control register signals to the out port
 -------------------------------------------------------------------------------
  INT_COUNT_PROCESS1: process (Clk)
  begin
    if (Clk'event and Clk = '1') then
      if (Rst = RESET_ACTIVE) then
        count <= (others => '1');
      elsif (Ld = '1') then
        count <= Load_in;
      elsif (En = '1' and zero_i = '0') then
          count <= count - 1;
      else
          null;
      end if;
    end if;
  end process INT_COUNT_PROCESS1;    
  
  INT_COUNT_PROCESS2: process (Clk)
  begin

    if (Clk'event and Clk = '1') then
      if (Rst = RESET_ACTIVE) then
        zero_i <= '1';
      else
        if (count = "00001") then
        zero_i <= '1';
        else
        zero_i <= '0';
        end if;
      end if;
    end if;
  end process INT_COUNT_PROCESS2;
  
  Zero <= zero_i;

end implementation;
